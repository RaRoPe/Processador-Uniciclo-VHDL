-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- ***************************************************************************
-- This file contains a Vhdl test bench template that is freely editable to   
-- suit user's needs .Comments are provided in each section to help the user  
-- fill out necessary details.                                                
-- ***************************************************************************
-- Generated on "02/06/2017 11:00:11"
                                                            
-- Vhdl Test Bench template for design  :  ANDBne
-- 
-- Simulation tool : ModelSim-Altera (VHDL)
-- 

LIBRARY ieee;                                               
USE ieee.std_logic_1164.all;                                

ENTITY ANDBne_tb IS
END ANDBne_tb;
ARCHITECTURE ANDBne_arch OF ANDBne_tb IS
-- constants                                                 
-- signals                                                   
SIGNAL andBne_out : STD_LOGIC;
SIGNAL bneControl : STD_LOGIC;
SIGNAL zeroULABne : STD_LOGIC;
COMPONENT ANDBne
	PORT (
	andBne_out : OUT STD_LOGIC;
	bneControl : IN STD_LOGIC;
	zeroULABne : IN STD_LOGIC
	);
END COMPONENT;
BEGIN
	i1 : ANDBne
	PORT MAP (
-- list connections between master ports and signals
	andBne_out => andBne_out,
	bneControl => bneControl,
	zeroULABne => zeroULABne
	);
init : PROCESS (bneControl, zeroULABne)
-- variable declarations                                     
BEGIN                                                        
        -- code that executes only once                      

END PROCESS init;                                           
always : PROCESS (bneControl, zeroULABne)
-- optional sensitivity list                                  
-- (        )                                                 
-- variable declarations                                      
BEGIN                                                         
        -- code executes for every event on sensitivity list  
		  bneControl <= '1';
		  zeroULABne <= '1';

END PROCESS always;                                          
END ANDBne_arch;
