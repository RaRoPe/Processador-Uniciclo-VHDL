-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- ***************************************************************************
-- This file contains a Vhdl test bench template that is freely editable to   
-- suit user's needs .Comments are provided in each section to help the user  
-- fill out necessary details.                                                
-- ***************************************************************************
-- Generated on "02/06/2017 03:17:52"
                                                            
-- Vhdl Test Bench template for design  :  pc
-- 
-- Simulation tool : ModelSim-Altera (VHDL)
-- 

LIBRARY ieee;                                               
USE ieee.std_logic_1164.all;                                

ENTITY pc_tb IS
END pc_tb;

ARCHITECTURE pc_arch OF pc_tb IS

	-- constants
	-- signals
	SIGNAL c_out : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL clk : STD_LOGIC;
	SIGNAL nextIns : STD_LOGIC_VECTOR(31 DOWNTO 0);

	COMPONENT pc
	
		PORT (
			c_out 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			clk 		: IN STD_LOGIC;
			nextIns 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
		
	END COMPONENT;

	BEGIN

		i1 : pc
		
		PORT MAP (
			-- list connections between master ports and signals
			c_out => c_out,
			clk => clk,
			nextIns => nextIns
		);
		
	init : PROCESS (clk, nextIns)
	-- variable declarations                                     
	
	BEGIN                                                        
			  -- code that executes only once                      
	
	END PROCESS init;                                           
	
	always : PROCESS (clk, nextIns)
	-- optional sensitivity list                                  
	-- (        )                                                 
	-- variable declarations                                      
	
	BEGIN                                                         
			  -- code executes for every event on sensitivity list  
			  clk <= '1';
			  nextIns <= "00000000000000000000000000000001";
	
	END PROCESS always;
	
END pc_arch;
