library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MODULO_SAIDA_INSTRUCTION is

	Port ( 
		SAIDA_INS_RS				: in STD_LOGIC_VECTOR (4 DOWNTO 0);
		SAIDA_INS_RT				: in STD_LOGIC_VECTOR (4 DOWNTO 0);
		SAIDA_INS_RD				: in STD_LOGIC_VECTOR (4 DOWNTO 0);
		SAIDA_INS_SHAMT			: in STD_LOGIC_VECTOR (4 DOWNTO 0);
		SAIDA_INS_FUNCT			: in STD_LOGIC_VECTOR (5 DOWNTO 0);
		SAIDA_INS_OPCODE			: in STD_LOGIC_VECTOR (5 DOWNTO 0);
		SAIDA_INS_IMM16			: in STD_LOGIC_VECTOR (15 DOWNTO 0);
		SAIDA_INS_IMM26			: in STD_LOGIC_VECTOR (25 DOWNTO 0);		
		
		-- V = VALOR DE SAIDA
		VSAIDA_INS_RS				: out STD_LOGIC_VECTOR (4 DOWNTO 0);
		VSAIDA_INS_RT				: out STD_LOGIC_VECTOR (4 DOWNTO 0);
		VSAIDA_INS_RD				: out STD_LOGIC_VECTOR (4 DOWNTO 0);
		VSAIDA_INS_SHAMT			: out STD_LOGIC_VECTOR (4 DOWNTO 0);
		VSAIDA_INS_FUNCT			: out STD_LOGIC_VECTOR (5 DOWNTO 0);
		VSAIDA_INS_OPCODE			: out STD_LOGIC_VECTOR (5 DOWNTO 0);
		VSAIDA_INS_IMM16			: out STD_LOGIC_VECTOR (15 DOWNTO 0);
		VSAIDA_INS_IMM26			: out STD_LOGIC_VECTOR (25 DOWNTO 0)
	);
	
end MODULO_SAIDA_INSTRUCTION;

architecture Behavioral of MODULO_SAIDA_INSTRUCTION is

begin
    
	VSAIDA_INS_RS			<= SAIDA_INS_RS;
	VSAIDA_INS_RT			<= SAIDA_INS_RT;
	VSAIDA_INS_RD			<= SAIDA_INS_RD;
	VSAIDA_INS_SHAMT		<= SAIDA_INS_SHAMT;
	VSAIDA_INS_FUNCT		<= SAIDA_INS_FUNCT;
	VSAIDA_INS_OPCODE		<= SAIDA_INS_OPCODE;
	VSAIDA_INS_IMM16		<= SAIDA_INS_IMM16;
	VSAIDA_INS_IMM26		<= SAIDA_INS_IMM26;
	 
end Behavioral;