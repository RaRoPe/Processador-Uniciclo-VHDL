library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity pc is

	Port ( 
		clk			: in  STD_LOGIC;
		nextIns		: in  STD_LOGIC_VECTOR (31 downto 0);
		c_out			: out STD_LOGIC_VECTOR (31 downto 0)
	);
	
end pc;

architecture Behavioral of pc is

begin
    c_out <= nextIns;
	 
end Behavioral;