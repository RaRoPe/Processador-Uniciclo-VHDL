library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MODULO_SAIDA is

	Port ( 
		SAIDA_PC				: in  STD_LOGIC_VECTOR (31 DOWNTO 0);
		SAIDA_MI				: in  STD_LOGIC_VECTOR (31 DOWNTO 0);
		SAIDA_MD				: in  STD_LOGIC_VECTOR (31 DOWNTO 0);
		SAIDA_BREG			: in  STD_LOGIC_VECTOR (31 DOWNTO 0);
		SAIDA_ULA			: in  STD_LOGIC_VECTOR (31 DOWNTO 0);
		SAIDA_SUMDESVIO	: in  STD_LOGIC_VECTOR (31 DOWNTO 0);
		SAIDA_SUMPC			: in  STD_LOGIC_VECTOR (31 DOWNTO 0);
		
		-- V = VALOR DE SAIDA
		VSAIDA_PC				: OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		VSAIDA_MI				: OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		VSAIDA_MD				: OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		VSAIDA_BREG				: OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		VSAIDA_ULA				: OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		VSAIDA_SUMDESVIO		: OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		VSAIDA_SUMPC			: OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	
end MODULO_SAIDA;

architecture Behavioral of MODULO_SAIDA is

begin
    
	VSAIDA_PC 				<= SAIDA_PC;
	VSAIDA_MI				<= SAIDA_MI;
	VSAIDA_MD				<= SAIDA_MD;
	VSAIDA_BREG				<= SAIDA_BREG;
	VSAIDA_ULA				<= SAIDA_ULA;
	VSAIDA_SUMDESVIO		<= SAIDA_SUMDESVIO;
	VSAIDA_SUMPC			<= SAIDA_SUMPC;
	 
end Behavioral;